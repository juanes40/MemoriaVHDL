library verilog;
use verilog.vl_types.all;
entity outputs_vlg_vec_tst is
end outputs_vlg_vec_tst;
